module rom(
    input wire clk,
    input wire [8:0] addr, // 9位地址可寻址512字
    output reg [31:0] data
);
    reg [31:0] mem [0:175];
    integer i;
    initial begin
        // 先全部清零
        for (i = 0; i < 176; i = i + 1) mem[i] = 32'b0;
        // jump.coe共44组，每组4个地址，原coe第n个值放到mem[n*4]
        mem[0]   = 32'h0100013c;
        mem[4]   = 32'h10000008;
        mem[8]   = 32'h00000000;
        mem[12]  = 32'h00000000;
        mem[16]  = 32'h00000000;
        mem[20]  = 32'h00000000;
        mem[24]  = 32'h00000000;
        mem[28]  = 32'h00000000;
        mem[32]  = 32'h1800000c;
        mem[36]  = 32'h0300013c;
        mem[40]  = 32'h00000000;
        mem[44]  = 32'h00000000;
        mem[48]  = 32'h00000000;
        mem[52]  = 32'h00000000;
        mem[56]  = 32'h00000000;
        mem[60]  = 32'h00000000;
        mem[64]  = 32'h20000234;
        mem[68]  = 32'h08004000;
        mem[72]  = 32'h0200013c;
        mem[76]  = 32'h00000000;
        mem[80]  = 32'h00000000;
        mem[84]  = 32'h00000000;
        mem[88]  = 32'h00000000;
        mem[92]  = 32'h00000000;
        mem[96]  = 32'h0f002214;
        mem[100] = 32'h0400013c;
        mem[104] = 32'h00000000;
        mem[108] = 32'h00000000;
        mem[112] = 32'h00000000;
        mem[116] = 32'h00000000;
        mem[120] = 32'h00000000;
        mem[124] = 32'h00000000;
        mem[128] = 32'h0600013c;
        mem[132] = 32'h21000008;
        mem[136] = 32'h00000000;
        mem[140] = 32'h00000000;
        mem[144] = 32'h00000000;
        mem[148] = 32'h00000000;
        mem[152] = 32'h00000000;
        mem[156] = 32'h00000000;
        mem[160] = 32'h0500013c;
        mem[164] = 32'h0500023c;
        mem[168] = 32'hf5ff2210;
        mem[172] = 32'h00000000;
    end
    reg [8:0] addr_r;
    always @(posedge clk) begin
        addr_r = addr;
        data = mem[addr_r];
    end
endmodule
