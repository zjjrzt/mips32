module rom(
    input wire clk,
    input wire [7:0] addr, // 9位地址可寻址512字
    output reg [31:0] data
);
    reg [31:0] mem [0:202]; // 203个值
    integer i;
    initial begin
        // 先全部清零
        for (i = 0; i < 203; i = i + 1) mem[i] = 32'b0;
        mem[0] = 32'h00608640;
        mem[1] = 32'h00688040;
        mem[2] = 32'h00010134;
        mem[3] = 32'h000001ac;
        mem[4] = 32'h00020134;
        mem[5] = 32'h0c000000;
        mem[6] = 32'h0000018c;
        mem[7] = 32'hffff023c;
        mem[8] = 32'h0080033c;
        mem[9] = 32'h20204300;
        mem[10] = 32'h00000000;
        mem[11] = 32'h00000000;
        mem[12] = 32'h00000000;
        mem[13] = 32'h00000000;
        mem[14] = 32'h00000000;
        mem[15] = 32'h00000000;
        mem[16] = 32'h00000000;
        mem[17] = 32'h00000000;
        mem[18] = 32'h00000000;
        mem[19] = 32'h00000000;
        mem[20] = 32'h4d000008;
        mem[21] = 32'h00000000;
        mem[22] = 32'h00000000;
        mem[23] = 32'h00000000;
        mem[24] = 32'h00000000;
        mem[25] = 32'h00000000;
        mem[26] = 32'h00000000;
        mem[27] = 32'h00000000;
        mem[28] = 32'h00000000;
        mem[29] = 32'h00000000;
        mem[30] = 32'h00000000;
        mem[31] = 32'h00000000;
        mem[32] = 32'h00000000;
        mem[33] = 32'h00000000;
        mem[34] = 32'h00000000;
        mem[35] = 32'h00000000;
        mem[36] = 32'h00000000;
        mem[37] = 32'h00000000;
        mem[38] = 32'h00000000;
        mem[39] = 32'h00000000;
        mem[40] = 32'h00000000;
        mem[41] = 32'h00000000;
        mem[42] = 32'h00000000;
        mem[43] = 32'h00000000;
        mem[44] = 32'h00000000;
        mem[45] = 32'h00000000;
        mem[46] = 32'h00000000;
        mem[47] = 32'h00000000;
        mem[48] = 32'h00000000;
        mem[49] = 32'h00000000;
        mem[50] = 32'h00000000;
        mem[51] = 32'h00000000;
        mem[52] = 32'h00000000;
        mem[53] = 32'h00000000;
        mem[54] = 32'h00000000;
        mem[55] = 32'h00000000;
        mem[56] = 32'h00000000;
        mem[57] = 32'h00000000;
        mem[58] = 32'h00000000;
        mem[59] = 32'h00000000;
        mem[60] = 32'h00000000;
        mem[61] = 32'h00000000;
        mem[62] = 32'h00000000;
        mem[63] = 32'h00000000;
        mem[64] = 32'h00680540;
        mem[65] = 32'h20000634;
        mem[66] = 32'h7d00a610;
        mem[67] = 32'h00000000;
        mem[68] = 32'h00680540;
        mem[69] = 32'h30000634;
        mem[70] = 32'h7900a610;
        mem[71] = 32'h00000000;
        mem[72] = 32'h4a000008;
        mem[73] = 32'h00000000;
        mem[74] = 32'hffff0734;
        mem[75] = 32'h4e000008;
        mem[76] = 32'h00000000;
        mem[77] = 32'h20204100;
        mem[78] = 32'h4e000008;
        mem[79] = 32'h00000000;
        mem[80] = 32'h00000000;
        mem[81] = 32'h00000000;
        mem[82] = 32'h00000000;
        mem[83] = 32'h00000000;
        mem[84] = 32'h00000000;
        mem[85] = 32'h00000000;
        mem[86] = 32'h00000000;
        mem[87] = 32'h00000000;
        mem[88] = 32'h00000000;
        mem[89] = 32'h00000000;
        mem[90] = 32'h00000000;
        mem[91] = 32'h00000000;
        mem[92] = 32'h00000000;
        mem[93] = 32'h00000000;
        mem[94] = 32'h00000000;
        mem[95] = 32'h00000000;
        mem[96] = 32'h00000000;
        mem[97] = 32'h00000000;
        mem[98] = 32'h00000000;
        mem[99] = 32'h00000000;
        mem[100] = 32'h00000000;
        mem[101] = 32'h00000000;
        mem[102] = 32'h00000000;
        mem[103] = 32'h00000000;
        mem[104] = 32'h00000000;
        mem[105] = 32'h00000000;
        mem[106] = 32'h00000000;
        mem[107] = 32'h00000000;
        mem[108] = 32'h00000000;
        mem[109] = 32'h00000000;
        mem[110] = 32'h00000000;
        mem[111] = 32'h00000000;
        mem[112] = 32'h00000000;
        mem[113] = 32'h00000000;
        mem[114] = 32'h00000000;
        mem[115] = 32'h00000000;
        mem[116] = 32'h00000000;
        mem[117] = 32'h00000000;
        mem[118] = 32'h00000000;
        mem[119] = 32'h00000000;
        mem[120] = 32'h00000000;
        mem[121] = 32'h00000000;
        mem[122] = 32'h00000000;
        mem[123] = 32'h00000000;
        mem[124] = 32'h00000000;
        mem[125] = 32'h00000000;
        mem[126] = 32'h00000000;
        mem[127] = 32'h00000000;
        mem[128] = 32'h00000000;
        mem[129] = 32'h00000000;
        mem[130] = 32'h00000000;
        mem[131] = 32'h00000000;
        mem[132] = 32'h00000000;
        mem[133] = 32'h00000000;
        mem[134] = 32'h00000000;
        mem[135] = 32'h00000000;
        mem[136] = 32'h00000000;
        mem[137] = 32'h00000000;
        mem[138] = 32'h00000000;
        mem[139] = 32'h00000000;
        mem[140] = 32'h00000000;
        mem[141] = 32'h00000000;
        mem[142] = 32'h00000000;
        mem[143] = 32'h00000000;
        mem[144] = 32'h00000000;
        mem[145] = 32'h00000000;
        mem[146] = 32'h00000000;
        mem[147] = 32'h00000000;
        mem[148] = 32'h00000000;
        mem[149] = 32'h00000000;
        mem[150] = 32'h00000000;
        mem[151] = 32'h00000000;
        mem[152] = 32'h00000000;
        mem[153] = 32'h00000000;
        mem[154] = 32'h00000000;
        mem[155] = 32'h00000000;
        mem[156] = 32'h00000000;
        mem[157] = 32'h00000000;
        mem[158] = 32'h00000000;
        mem[159] = 32'h00000000;
        mem[160] = 32'h00000000;
        mem[161] = 32'h00000000;
        mem[162] = 32'h00000000;
        mem[163] = 32'h00000000;
        mem[164] = 32'h00000000;
        mem[165] = 32'h00000000;
        mem[166] = 32'h00000000;
        mem[167] = 32'h00000000;
        mem[168] = 32'h00000000;
        mem[169] = 32'h00000000;
        mem[170] = 32'h00000000;
        mem[171] = 32'h00000000;
        mem[172] = 32'h00000000;
        mem[173] = 32'h00000000;
        mem[174] = 32'h00000000;
        mem[175] = 32'h00000000;
        mem[176] = 32'h00000000;
        mem[177] = 32'h00000000;
        mem[178] = 32'h00000000;
        mem[179] = 32'h00000000;
        mem[180] = 32'h00000000;
        mem[181] = 32'h00000000;
        mem[182] = 32'h00000000;
        mem[183] = 32'h00000000;
        mem[184] = 32'h00000000;
        mem[185] = 32'h00000000;
        mem[186] = 32'h00000000;
        mem[187] = 32'h00000000;
        mem[188] = 32'h00000000;
        mem[189] = 32'h00000000;
        mem[190] = 32'h00000000;
        mem[191] = 32'h00000000;
        mem[192] = 32'h0100e724;
        mem[193] = 32'h00700940;
        mem[194] = 32'h04000834;
        mem[195] = 32'h20482801;
        mem[196] = 32'h00708940;
        mem[197] = 32'h00000000;
        mem[198] = 32'h18000042;
        mem[199] = 32'h00000000;
        mem[200] = 32'h00000000;
        mem[201] = 32'h00000000;
        mem[202] = 32'h00000000;
    end
    reg [8:0] addr_r;
    always @(posedge clk) begin
        addr_r = addr;
        data = mem[addr_r];
    end
endmodule
