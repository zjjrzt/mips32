//取指/译码寄存器模块

module ifid_reg(
    input wire clk,
    input wire rst_n,
    input wire [31:0] if_pc,        //取指阶段的pc值
    output reg [31:0] id_pc        //译码阶段的pc值
);


    always @(posedge clk or negedge rst_n) begin
        if(!rst_n) begin
            id_pc <= 32'h0000_3000;
        end
        else begin
            id_pc <= if_pc;
        end
    end

endmodule